��  CCircuit��  CSerializeHack           ��  CPart              ��� 	 CResistor��  CValue  � i� w    200           i@      �?   �� 	 CTerminal  � P� e         ������@�'m�?  �  � |� �      	 -�ZL��?�'m��    � d� |         ��      ��  CBattery
�  k���    3.7V(    ������@      �? V �  �p��         ������@�Iu���ɿ  �  ����                �Iu����?    ����         ��      ��  CNPN��  CDummyValue  ��    100hFE            Y@      �? hFE �  p�       	 b���^�?T^����?  �  � �� �        -�ZL��?�'m�?  �  ��                 �<u���ɿ    � ��         ��      ��  CDiode�  HTIi        b���^�?�A+�+�  �  H(I=         ������@�A+�+�=    <<TT        ��      ��  CMotorEM�  0E         ������@ ������?  �  \q        b���^�? �����ǿ  �� 	 CMechTerm�Ǭ�G���^�#`Z��      �<                  @!E     	 �Ǭ�G��      �<    D\     !   ��      bK�6�>�Ǭ�G���^	����fF�h��!��Ǭ�G���^	����              ���  CWire  (I)      &�  � ()      &�  � (� Q       &�  ���       &�  H(�)      &�  �(�q       &�  hIi      &�  pq      &�  hq       &�  (1                     �                             )      ,    *  "       *   -  '  ! 0 ! " " . $ $   0 + ) ' (     , +  /   / - . ( !           �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 