��  CCircuit��  CSerializeHack           ��  CPart              ���  CDiode�� 	 CTerminal  $9        {�;)�?�0]����  
�  �          ������@�0]����=    $$        ��      ��  CBattery��  CValue  39[G    3.7V(    ������@      �? V 
�  h i5         ������@0�'j:�ǿ  
�  hLia                 0�'j:��?    \4tL         ��      ��  CMotorEM
�  � � �          ������@�K�i:��?  
�  � $� 9        {�;)�?�K�i:�ǿ  �� 	 CMechTerm>�1+�����qk4+��      �<                  �      	 >�1+����      �<    � � $        ��      bK�6�>>�1+������E����bT42�!�>�1+������E������  S q{     5V(          @      �? V 
�  � X� m       	       @���E^q�  
�  � �� �                ���E^q?    | l� �         ��      �� 	 CResistor�  � F� T    1k        @�@      �?k  
�  � X� Y        �(p�Q�?���E^q�  
�  � X� Y              @���E^q?    � T� \         ��      ��  CNPN��  CDummyValue  � H� H    100hFE            Y@      �? hFE 
�  � 8� M       	 {�;)�?v�'j:��?  
�  � X� Y      	 �(p�Q�?���E^q?  
�  � d� y                 ��T�*;ȿ    � L� d     &    ��                    ���  CWire  � i�       *�  � 89      *�  � � �       *�  � �i�       *�  � �� �       *�  � x� �        *�  h`i�        *�  h� i!                     �                              ,  +   2    1  -    &      !    /     ' !  ! & , & '   ' ( ( 0 - 2     / 1  0 ( .  . +            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 