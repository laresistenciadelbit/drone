��  CCircuit��  CSerializeHack           ��  CPart              ���  CBulb�� 	 CTerminal  � �� �               @�Q���?  
�  � ��                ��Q��롿    � �� �        ��      ��  CBattery��  CValue  C k     3.5V(          @      �? V 
�  x �y �               @�Q��뱿  
�  x y )               ��Q���?    l ��          ��      �
�  � �� �               @�Q���?  
�  � ��                ��Q��롿    � �� �        ��      ��  CDiode
�  ����                Ɯ�C�  
�  ����               @Ɯ�C�=    ����        ��      ��  ���    3.5V(          @      �? V 
�   �!�               @+On/���  
�   !                +On/��@    �,         ��      �� 	 CResistor�  ����    1.35     �������?      �?   
�  ����               @�Kh/��@  
�  ����                �Kh/���    ����     !    ��      ��  CNPN��  CExplode              �p ͦs@       @ A��  CDummyValue   ( (    100hFE            Y@      �? hFE 
�   -       	 ������@         
�  �8�9      	 ffffff
@         
�   DY       	                    �,D     )    ��      ��  �&�4    1         �?      �?   
�  �8�9        ffffff
@          
�  �8�9        ffffff
@            �4�<    .    ��      ��  cQ�_    3.3V(    ffffff
@      �? V 
�  �8�M       	 ffffff
@          
�  �d�y                            �L�d     2    ��      ��  CMotorEM
�   � �          ������@����ѣ�  
�           ������@����ѣ<  �� 	 CMechTermNY6�=        p��xs"�                  � �      	 NY6�=p��xs"�    ��      6   ��      bK�6�>NY6�=�4(D�(�     �v�NY6�=�4(D�(���  Ck'    3.7V(    ������@      �? V 
�  x y         ������@��� �ѣ<  
�  x,yA                 ��� �ѣ�    l�,     <    ��      �
�  ()        ������@�i�c�A;  
�  (� )�          ������@�i�c�A�    � 4    ?    ��      ��  {	�    1.35     �������?      �?   
�  �� �         ����@����L9�?  
�  ��1        	!�m��
@����L9п    ��     C    ��      #�'�  �@�@    100hFE            Y@      �? hFE 
�  �0�E       	 	!�m��
@M���L9�?  
�  xP�Q     	 	 !��{�?{'��9�d?  
�  �\�q          �̰Ծ�af�bп    �D�\     G    ��      ��  H>hL    1k        @�@      �?k  
�  dPyQ     	   !��{�?>'��9�d�  
�  8PMQ     
   ��L�cf
@>'��9�d?    LLdT    L    ��      ��  i+w    3.3V(    ffffff
@      �? V 
�  8P9e      
 	 ��L�cf
@>'��9�d�  
�  8|9�         �̰Ծ��9�d?    ,dD|     P    ��      ��  �1?    3.7V(    ������@      �? V 
�  -         ����@����L9п  
�  DY          �̰Ծz���L9�?    ,$D     T    ��      �
�  ��1        	!�m��
@R�T�Vв�  
�  �� �         ����@R�T�Vв=    ��    W    ��      �
�  $9        ��~��v?�`���d�  
�  �          ��a��@�`���d�=    $$    Z    ��      ��  39[G    3.7V(    ������@      �? V 
�  h i5         ��a��@���'�#ȿ  
�  hLia         P���$G?�,�'�#�?    \4tL     ^    ��      4�
�  � � �          ��a��@�hV'�#�?  
�  � $� 9        ��~��v?�hV'�#ȿ  8���[P�	� ����      Լ                  �      	 ��[P�	�      Լ    � � $     a   ��      bK�6�>��[P�	�����[8�4�1_�!���[P�	�����[8���  S q{     3.3V(    ffffff
@      �? V 
�  � X� m       	 {�.��g
@%l ͦs�  
�  � �� �         P���$G?@o ͦs@    | l� �     f    ��      ��  � F� T    1         �?      �?   
�  � X� Y        ��8����?|p ͦs�  
�  � X� Y        {�.��g
@|p ͦs@    � T� \    j    ��      #�'�  � H� H    100hFE            Y@      �? hFE 
�  � 8� M       	 ��~��v? �'�#�?  
�  � X� Y      	 ��8����?ip ͦs@  
�  � d� y         P���$G?2�����    � L� d     n    ��                    ���  CWire  x (� )      r�  � � )       r�  � �       r�  � �� �      r�  x �� �      r�  x �y �       r�  ����      r�  ����      r�  ���       r�  �!      r�  � i�       r�  ��!�      r�   �!�       r�  ����      r�  x� y       r�  x@yy        r�   Xy        r�  �xy       r�   xyy       r�   � )�       r�   )      r�  (� y�       r�  �� ��       r�  �        r�  X�       r�  �p��       r�  8���      r�  ���      r�  �0�1      r�  �� �       r�  � 89      r�  � � �       r�  � �i�      r�  � �� �      r�  � x� �       r�  h`i�       r�  h� i!                     �                             v    u  x    s  w    u   y  ~       | ! � ! " " z ) � ) * . * + + � . . * / 2 / 2 / 2 3 3 � 6 � 6 7 7 ) 9 9   < � < = = � ? ? � @ � @ C � C D D G G � G H L H I I � L L H M P M P M P Q Q � T � T U U � W W � X � X Z Z � [ } [ ^ � ^ _ _ � a � a b b n c c   f k f g g � j j o k f k n � n o j o p p �  t  s t    x v w  z  " { y | {  � � �  ~  !  � < = � + � 3 � � � 6 @ 7 ? � � C X � T U � I � Q � � � D W � � b Z a [ � � g � p � _ � } ^   0        �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 